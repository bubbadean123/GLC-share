module instruction_decoder(instruction,r_zero, load_a, load_b, load_r, jump_up, jump_dowm, b_immediate, ivalue );

endmodule